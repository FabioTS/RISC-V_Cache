library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.constants.all;

entity cache is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity cache;

architecture RTL of cache is
	
begin

end architecture RTL;
